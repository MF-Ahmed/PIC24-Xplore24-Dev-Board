** Profile: "SCHEMATIC1-Bias"  [ C:\My Documents\z02-schematic1-bias.sim ] 

** Creating circuit file "z02-schematic1-bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.OP
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\Z02-SCHEMATIC1.net" 


.END
